module exu (
    
);
    
    
endmodule