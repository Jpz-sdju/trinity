module issuequeue (
    
);
    
endmodule