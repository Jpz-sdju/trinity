`include "defines.sv"
module mshr_entry (
    input wire                clock,          // Clock signal
    input wire                reset_n,        // Active low reset
    input wire                install_valid,
    input wire [`PADDR_RANGE] install_paddr


);

endmodule
