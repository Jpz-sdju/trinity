module storeunit (
    
);
    
endmodule